`ifndef __AUDIO_DEFS_VH__
`define __AUDIO_DEFS_VH__

localparam int DFX_REG_CTRL           = 0;
localparam int STEREO                 = 1;
localparam int AUDIO_WIDTH            = 24;

`endif // AUDIO_DEFS_VH
