`ifndef __LP_DEFS_VH__
`define __LP_DEFS_VH__

`endif // __LP_DEFS_VH__
