`ifndef __DSD_DEFS_VH__
`define __DSD_DEFS_VH__

`define AUDIO_IN = 24;
`define NCOEFFS = 500;
`define COEFF_W = 32;
`define INITIAL_COEFFS = "dsd_coeff_32.hex";

`endif // DSD_DEFS_VH
