// ------------------------------------------------------------------------
// Filename:       llac_audio_system_top.sv
//
// Project:        LLAC, intelligent hardware scheduler targeting common
// audio signal chains.
//
// For more information see the repository:
// https://github.com/topologicalhurt/Thesis
//
// Purpose:        N/A
//
// Author: topologicalhurt csin0659@uni.sydney.edu.au
//
// ------------------------------------------------------------------------
// Copyright (C) 2025, LLAC project LLC
//
// This file is a part of the RTL module
// It is intended to be used as part of the Out design where a README.md
// detailing the design should exist, conforming to the details provided
// under docs/CONTRIBUTING.md. The Out module is covered by the GPL 3.0
// License (see below.)
//
// The design is NOT COVERED UNDER ANY WARRANTY.
//
// LICENSE:     GNU GENERAL PUBLIC LICENSE Version 3, 29 June 2007
// As defined by GNU GPL 3.0 https://www.gnu.org/licenses/gpl-3.0.html
//
// A copy of this license is included at the root directory. It should've
// been provided to you
// Otherwise please consult:
// https://github.com/topologicalhurt/Thesis/blob/main/LICENSE
// ------------------------------------------------------------------------


module llac_audio_system_top #(
    parameter int NUM_CORES = 4,
    parameter int AUDIO_WIDTH = 24,
    parameter int AXI_ADDR_WIDTH = 32,
    parameter int AXI_DATA_WIDTH = 64,
    parameter int AXI_ID_WIDTH = 6
) (
    // Clocks and reset
    input  logic        clk_100mhz,   // 100MHz system clock from PYNQ-Z2
    input  logic        clk_audio,    // Audio clock (typically 24.576MHz for 48kHz)
    input  logic        resetn,       // Active low reset

    // Audio core bus signals
    input logic [NUM_CORES-1:0]       core_pause,
    input logic [NUM_CORES-1:0]       core_stop,
    input logic [NUM_CORES-1:0]       core_resume,
    input logic [NUM_CORES-1:0]       core_status,
    input logic [NUM_CORES-1:0]       core_interrupt,

    // AXI4 memory interface for DRAM
    // Write Address Channel
    output logic [AXI_ID_WIDTH-1:0]        m_axi_awid,
    output logic [AXI_ADDR_WIDTH-1:0]      m_axi_awaddr,
    output logic [7:0]                     m_axi_awlen,
    output logic [2:0]                     m_axi_awsize,
    output logic [1:0]                     m_axi_awburst,
    output logic                           m_axi_awlock,
    output logic [3:0]                     m_axi_awcache,
    output logic [2:0]                     m_axi_awprot,
    output logic [3:0]                     m_axi_awqos,
    output logic                           m_axi_awvalid,
    input  logic                           m_axi_awready,

    // Write Data Channel
    output logic [AXI_DATA_WIDTH-1:0]      m_axi_wdata,
    output logic [AXI_DATA_WIDTH/8-1:0]    m_axi_wstrb,
    output logic                           m_axi_wlast,
    output logic                           m_axi_wvalid,
    input  logic                           m_axi_wready,

    // Write Response Channel
    input  logic [AXI_ID_WIDTH-1:0]        m_axi_bid,
    input  logic [1:0]                     m_axi_bresp,
    input  logic                           m_axi_bvalid,
    output logic                           m_axi_bready,

    // Read Address Channel
    output logic [AXI_ID_WIDTH-1:0]        m_axi_arid,
    output logic [AXI_ADDR_WIDTH-1:0]      m_axi_araddr,
    output logic [7:0]                     m_axi_arlen,
    output logic [2:0]                     m_axi_arsize,
    output logic [1:0]                     m_axi_arburst,
    output logic                           m_axi_arlock,
    output logic [3:0]                     m_axi_arcache,
    output logic [2:0]                     m_axi_arprot,
    output logic [3:0]                     m_axi_arqos,
    output logic                           m_axi_arvalid,
    input  logic                           m_axi_arready,

    // Read Data Channel
    input  logic [AXI_ID_WIDTH-1:0]        m_axi_rid,
    input  logic [AXI_DATA_WIDTH-1:0]      m_axi_rdata,
    input  logic [1:0]                     m_axi_rresp,
    input  logic                           m_axi_rlast,
    input  logic                           m_axi_rvalid,
    output logic                           m_axi_rready,

    // AXI4-Lite slave interface for control
    input  logic [AXI_ADDR_WIDTH-1:0]      s_axil_awaddr,
    input  logic                           s_axil_awvalid,
    output logic                           s_axil_awready,

    input  logic [31:0]                    s_axil_wdata,
    input  logic [3:0]                     s_axil_wstrb,
    input  logic                           s_axil_wvalid,
    output logic                           s_axil_wready,

    output logic [1:0]                     s_axil_bresp,
    output logic                           s_axil_bvalid,
    input  logic                           s_axil_bready,

    input  logic [AXI_ADDR_WIDTH-1:0]      s_axil_araddr,
    input  logic                           s_axil_arvalid,
    output logic                           s_axil_arready,

    output logic [31:0]                    s_axil_rdata,
    output logic [1:0]                     s_axil_rresp,
    output logic                           s_axil_rvalid,
    input  logic                           s_axil_rready,

    // Interrupt
    output logic                           irq_out,

    // I2S interface signals
    output logic                           i2s_mclk,      // Master clock (optional)
    output logic                           i2s_bclk,      // Bit clock
    output logic                           i2s_lrclk,     // Left/Right clock (Word Select)
    input  logic                           i2s_sdata_in,  // Serial data input from ADC
    output logic                           i2s_sdata_out, // Serial data output to DAC

    // I2C control interface for codec configuration
    inout  wire                            i2c_scl,
    inout  wire                            i2c_sda,

    // Debug/Status LEDs
    output logic [3:0]                     leds
);
    // Local parameters
    localparam int CORE_ID_WIDTH = $clog2(NUM_CORES);

    // Audio data signals
    logic [AUDIO_WIDTH-1:0]     audio_left_in;
    logic [AUDIO_WIDTH-1:0]     audio_right_in;
    logic [AUDIO_WIDTH-1:0]     audio_left_out;
    logic [AUDIO_WIDTH-1:0]     audio_right_out;
    logic                       audio_valid_in;
    logic                       audio_valid_out;
    logic                       audio_ready_in;
    logic                       audio_ready_out;

    // Fifo status
    logic                       fifo_overflow;
    logic                       fifo_underflow;
    logic [3:0]                 dac_status;

    // Generate master clock for audio codec (typically 256fs or 512fs)
    // Assuming clk_audio is already the correct frequency
    assign i2s_mclk = clk_audio;

    // Forward status to LEDs for debugging
    assign leds = dac_status;

    // Audio DAC Interface
    audio_dac_interface #(
        .AUDIO_DATA_WIDTH(AUDIO_WIDTH)
    ) dac_interface (
        .clk_100mhz(clk_100mhz),
        .resetn(resetn),
        .audio_clk(clk_audio),

        // Audio data input
        .audio_left_in(audio_left_out),
        .audio_right_in(audio_right_out),
        .audio_valid_in(audio_valid_out),
        .audio_ready_out(audio_ready_out),

        // I2S signals to codec
        .i2s_bclk(i2s_bclk),
        .i2s_lrclk(i2s_lrclk),
        .i2s_sdata(i2s_sdata_out),

        // I2C control interface
        .i2c_scl(i2c_scl),
        .i2c_sda(i2c_sda),

        // Status signals
        .fifo_overflow(fifo_overflow),
        .fifo_underflow(fifo_underflow),
        .status(dac_status)
    );

    // Audio input processor
    buf_audio_in #(
        .I2S_WIDTH(AUDIO_WIDTH),
        .NUM_AUDIO_CHANNELS(NUM_CORES)
    ) adc_interface (
        .sys_clk(clk_100mhz),
        .sys_rst(~resetn),

        // I2S Interface (from external ADC)
        .i2s_bclk(i2s_bclk),
        .i2s_lrclk(i2s_lrclk),
        .i2s_data(i2s_sdata_in),

        // Output valid signal
        .sample_valid(audio_valid_in)
    );

    // Main system interface for control and memory access
    llac_top_interface #(
        .NUM_CORES(NUM_CORES),
        .NUM_INTERRUPTS(8),
        .AXI_ID_WIDTH(AXI_ID_WIDTH),
        .AXI_ADDR_WIDTH(AXI_ADDR_WIDTH),
        .AXI_DATA_WIDTH(AXI_DATA_WIDTH)
    ) top_if (
        .clk(clk_100mhz),
        .resetn(resetn),

        // AXI4 Memory Interface
        .m_axi_awid(m_axi_awid),
        .m_axi_awaddr(m_axi_awaddr),
        .m_axi_awlen(m_axi_awlen),
        .m_axi_awsize(m_axi_awsize),
        .m_axi_awburst(m_axi_awburst),
        .m_axi_awlock(m_axi_awlock),
        .m_axi_awcache(m_axi_awcache),
        .m_axi_awprot(m_axi_awprot),
        .m_axi_awqos(m_axi_awqos),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awready(m_axi_awready),

        .m_axi_wdata(m_axi_wdata),
        .m_axi_wstrb(m_axi_wstrb),
        .m_axi_wlast(m_axi_wlast),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),

        .m_axi_bid(m_axi_bid),
        .m_axi_bresp(m_axi_bresp),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready),

        .m_axi_arid(m_axi_arid),
        .m_axi_araddr(m_axi_araddr),
        .m_axi_arlen(m_axi_arlen),
        .m_axi_arsize(m_axi_arsize),
        .m_axi_arburst(m_axi_arburst),
        .m_axi_arlock(m_axi_arlock),
        .m_axi_arcache(m_axi_arcache),
        .m_axi_arprot(m_axi_arprot),
        .m_axi_arqos(m_axi_arqos),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arready(m_axi_arready),

        .m_axi_rid(m_axi_rid),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rresp(m_axi_rresp),
        .m_axi_rlast(m_axi_rlast),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready),

        // AXI4-Lite Control Interface
        .s_axil_awaddr(s_axil_awaddr),
        .s_axil_awvalid(s_axil_awvalid),
        .s_axil_awready(s_axil_awready),

        .s_axil_wdata(s_axil_wdata),
        .s_axil_wstrb(s_axil_wstrb),
        .s_axil_wvalid(s_axil_wvalid),
        .s_axil_wready(s_axil_wready),

        .s_axil_bresp(s_axil_bresp),
        .s_axil_bvalid(s_axil_bvalid),
        .s_axil_bready(s_axil_bready),

        .s_axil_araddr(s_axil_araddr),
        .s_axil_arvalid(s_axil_arvalid),
        .s_axil_arready(s_axil_arready),

        .s_axil_rdata(s_axil_rdata),
        .s_axil_rresp(s_axil_rresp),
        .s_axil_rvalid(s_axil_rvalid),
        .s_axil_rready(s_axil_rready),

        // Interrupt
        .irq_out(irq_out),

        // Audio interface
        .audio_clk(clk_audio),
        .audio_rst(~resetn),

        // Core control
        .core_pause(core_pause),
        .core_stop(core_stop),
        .core_resume(core_resume),
        .core_status(core_status),
        .core_interrupt(core_interrupt)
    );

    // Audio processing cores
    // In a real implementation, these would be the dynamically reconfigurable audio cores
    // For simplicity, this example just has some placeholders

    // Passthrough
    always_ff @(posedge clk_100mhz or negedge resetn) begin
        if (!resetn) begin
            audio_left_out <= '0;
            audio_right_out <= '0;
            audio_valid_out <= 1'b0;
            core_status <= '0;
            core_interrupt <= '0;
        end else begin
            // Basic passthrough logic
            if (audio_valid_in && audio_ready_out) begin
                // Extract input from first audio channel
                // In real implementation, this would go through the ensemble cores
                audio_left_out <= audio_left_out[0];
                audio_right_out <= audio_right_out[0];
                audio_valid_out <= 1'b1;

                // Signal that core is active
                core_status[0] <= 1'b1;
            end else begin
                audio_valid_out <= 1'b0;
            end

            // Handle core control signals
            for (int i = 0; i < NUM_CORES; i++) begin
                if (core_pause[i]) begin
                    core_status[i] <= 1'b0;  // Mark as paused
                end
                if (core_stop[i]) begin
                    core_status[i] <= 1'b0;  // Mark as stopped
                    core_interrupt[i] <= 1'b1;  // Signal completion
                end
                if (core_resume[i]) begin
                    core_status[i] <= 1'b1;  // Mark as active
                    core_interrupt[i] <= 1'b0;  // Clear interrupt
                end
            end
        end
    end

endmodule : llac_audio_system_top
