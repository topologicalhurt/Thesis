`ifndef __SINC_DEFS_VH__
`define __SINC_DEFS_VH__

`define N_STAGES = 5 // Number of approximation stages (design accumulates as power of 2) I.e. 5 => 2^5 = 32
`define AUDIO_WIDTH = 24

`endif // __SINC_DEFS_VH__
