`ifndef CORE_CONSTS_SVH
`define CORE_CONSTS_SVH

`define PI_OVER_2         24'd1647099   // π/2 in Q2.22
`define PI                24'd3294198   // π   in Q2.22
`define THREE_PI_OVER_2   24'd4941297   // 3π/2 in Q2.22
`define TWO_PI            24'd6588396   // 2π in Q2.22 (optional)

`endif // CORE_CONSTS_SVH
