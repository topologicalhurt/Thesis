`ifndef __DSD_DEFS_VH__
`define __DSD_DEFS_VH__

localparam int NCOEFFS      = 500;
localparam int COEFF_W      = 32;
parameter      INITIAL_COEFFS = "dsd_coeff_32.hex";

`endif // DSD_DEFS_VH
