`ifndef __AUDIO_DEFS_VH__
`define __AUDIO_DEFS_VH__

// Audio buffer configuration parameters
localparam int DFX_REG_CTRL           = 0;
localparam int STEREO                 = True;
localparam int AUDIO_WIDTH            = 24;
localparam int BUFFER_DEPTH           = 4;

`endif // AUDIO_DEFS_VH
