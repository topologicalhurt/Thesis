`ifndef __AVG_IIR_TB_VH__
`define __AVG_IIR_TB_VH__

`endif // __AVG_IIR_TB_VH__
