`ifndef __HP_DEFS_VH__
`define __HP_DEFS_VH__

`endif // __HP_DEFS_VH__
