`ifndef __AVG_IIR_DEFS_VH__
`define __AVG_IIR_DEFS_VH__

`endif // __AVG_IIR_DEFS_VH__
