`ifndef __DSD_TB_VH__
`define __DSD_TB_VH__

`endif // __DSD_TB_VH__
